`ifndef __MUNOC_ROUTER_ID_H__
`define __MUNOC_ROUTER_ID_H__

`define ROUTER_ID_I_SYSTEM_ROUTER (0)

`endif