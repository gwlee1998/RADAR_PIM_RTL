`ifndef __USER_INFO_H__
`define __USER_INFO_H__



`endif