`ifndef __IROM_CAPACITY_H__
`define __IROM_CAPACITY_H__

`define IROM_CAPACITY 648

`endif