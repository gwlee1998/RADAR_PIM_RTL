wire [BW_USERNAME-1:0] username_string = `FORMAT_STRING("cau1_lab11");
wire [BW_GIT_NAME-1:0] home_git_name_string = `FORMAT_STRING("rvx_dev");
wire [BW_GIT_VERSION-1:0] home_git_version_string = `FORMAT_STRING("9b0c9d4");
wire [BW_GIT_VERSION-1:0] devkit_git_version_string = `FORMAT_STRING("509d0ef");
wire [BW_DATE-1:0] design_date_string = `FORMAT_STRING("2023-11-23 10:09");