`ifndef __PLATFORM_INFO_H__
`define __PLATFORM_INFO_H__

`include "memorymap_info.vh"
`include "hw_info.vh"
`include "ssw_info.vh"
`include "user_info.vh"


`endif